--------------------------------------------------
-- Project: Black-jack
-- File:  card_deck.vhd
-- Authors: Daiane Fraga, George Redivo
--------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_arith.all;
    use ieee.std_logic_unsigned.all;   

entity card_deck is
    Port ( 	
				clk : in  STD_LOGIC;
				rst : in  STD_LOGIC;
				card_out: out  STD_LOGIC_VECTOR(3 downto 0)
			);
end card_deck;

architecture card_deck of card_deck is

type card_bank is array(51 downto 0) of std_logic_vector(3 downto 0);

signal sig_card_out : std_logic_vector(3 downto 0);
signal card : card_bank;
signal counter : integer;

constant NUMBER_OF_CARDS : integer := 52;

begin
	-- Paste here the code generated by program shuffle
	card(0) <= "0010"; -- 2
	card(1) <= "0011"; -- 3
	card(2) <= "0101"; -- 5
	card(3) <= "0110"; -- 6
	card(4) <= "0110"; -- 6
	card(5) <= "1000"; -- 8
	card(6) <= "1010";
	card(7) <= "1100";
	card(8) <= "0011";
	card(9) <= "1001";
	card(10) <= "1101";
	card(11) <= "0111";
	card(12) <= "0010";
	card(13) <= "1010";
	card(14) <= "0111";
	card(15) <= "0111";
	card(16) <= "1011";
	card(17) <= "1101";
	card(18) <= "1001";
	card(19) <= "0010";
	card(20) <= "1100";
	card(21) <= "0001";
	card(22) <= "0101";
	card(23) <= "1010";
	card(24) <= "0110";
	card(25) <= "1010";
	card(26) <= "0001";
	card(27) <= "1011";
	card(28) <= "1001";
	card(29) <= "0100";
	card(30) <= "0010";
	card(31) <= "0100";
	card(32) <= "1000";
	card(33) <= "0001";
	card(34) <= "0001";
	card(35) <= "0101";
	card(36) <= "1001";
	card(37) <= "1101";
	card(38) <= "1011";
	card(39) <= "0011";
	card(40) <= "1000";
	card(41) <= "0110";
	card(42) <= "1100";
	card(43) <= "0111";
	card(44) <= "1101";
	card(45) <= "1011";
	card(46) <= "0100";
	card(47) <= "0100";
	card(48) <= "1100";
	card(49) <= "1000";
	card(50) <= "0101";
	card(51) <= "0011";
	-- end of paste

  card_out <= sig_card_out;
  
	process (clk, rst)
	begin
		if (clk'event and clk = '1') then
			if rst = '1' then
				counter <= 0;
			elsif (counter >= 0 and counter < NUMBER_OF_CARDS) then
				sig_card_out <= card(counter);
				counter <= counter + 1;
			else
				counter <= 0;
        -- This causes invalid index on the vector...
				--sig_card_out <= card(counter);
			end if;
		end if;
	end process;

end card_deck;

