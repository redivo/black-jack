--------------------------------------------------
-- Project: Black-jack
-- File:  card_deck.vhd
-- Authors: Daiane Fraga, George Redivo
--------------------------------------------------
library ieee;
    use ieee.std_logic_1164.all;
    use ieee.std_logic_arith.all;
    use ieee.std_logic_unsigned.all;   


entity card_deck is
    Port ( 	
				clk : in  STD_LOGIC;
				rst : in  STD_LOGIC;
				card_out: out  STD_LOGIC_VECTOR(3 downto 0)
			);
end card_deck;

architecture card_deck of card_deck is

type card_bank is array(51 downto 0) of std_logic_vector(3 downto 0);

signal sig_card_out : std_logic_vector(3 downto 0);
signal card : card_bank;
signal counter : integer;

constant NUMBER_OF_CARDS : integer := 52;

begin
	-- Paste here the code generated by program shuffle

	-- end of paste

	process (clk, rst)
	begin
		if (clk'event and clk = '1') then
			if counter < NUMBER_OF_CARDS then
				sig_card_out <= card(counter);
				counter <= counter + 1;
			else
				counter <= 0;
				sig_card_out <= card(counter);
			end if;
		end if;
	end process;

end card_deck;

