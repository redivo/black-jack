----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Daiane Fraga, George Pinto
-- 
-- Create Date:    18:28:52 05/19/2013 
-- Design Name: 
-- Module Name:    card deck
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: Module to load the cards
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity card_deck is
    Port ( clk : in  STD_LOGIC;
           card_out: out  STD_LOGIC_VECTOR(3 downto 0));
end card_deck;

architecture card_deck of card_deck is

type card_bank is array(51 downto 0) of std_logic_vector(3 downto 0);

signal sig_card_out : std_logic_vector(3 downto 0);
signal card : card_bank;
signal counter : integer;

constant NUMBER_OF_CARDS : integer := 52;

begin
	-- Paste here the code generated by program shuffle

	-- end of paste

	process (clk, rst)
	begin
		if (clk'event and clk = '1') then
			if counter < NUMBER_OF_CARDS then
				sig_card_out <= card(counter);
				counter <= counter + 1;
			else
				counter = 0;
				sig_card_out <= card(counter);
			end if;
		end if;
	end process;

end card_deck;

